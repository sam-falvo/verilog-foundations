module queue(
);

endmodule

